library IEEE;
use IEEE.Std_Logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity decod is port (
	A: in std_logic_vector (3 downto 0);
);

architecture decod_arch of decod is begin

end decod_arch;