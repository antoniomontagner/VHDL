library IEEE;
use IEEE.std_logic_1164.all

entity tb_contador is 
end tb_contador;

architecture bvh of tb_contador is

    signal clk : std_logic;
    signal q: unsigned (3 downto 0);

begin


end bvh ; 